//------------------------------------------------------------------------------
//	Module:		LevelToPulse
//	Desc:			This module provides a 1-cycle output based on a push button
//					raw input source.
//	Params:		This module is not parameterized.
//	Inputs:		See Lab2 document
//	Outputs:		See Lab2 document
//
//	Author:     LUCAS OLIVEIRA SILVA
//				LUCAS HENRIQUE COSTA ARAUJO
//------------------------------------------------------------------------------
module	LevelToPulse(
			//------------------------------------------------------------------
			//	Clock & Reset Inputs
			//------------------------------------------------------------------
			 Clock,
			 Reset,
			//------------------------------------------------------------------
			

			//------------------------------------------------------------------
			//	Inputs
			//------------------------------------------------------------------
			 Level,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Outputs
			//------------------------------------------------------------------
			 Pulse 
			//------------------------------------------------------------------
	);

	
	//--------------------------------------------------------------------------
	//	Clock & Reset Inputs
	//--------------------------------------------------------------------------
	input					Clock;	// System clock
	input					Reset;	// System reset
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Inputs
	//--------------------------------------------------------------------------
	input					Level;
	//--------------------------------------------------------------------------


	//--------------------------------------------------------------------------
	//	Outputs
	//--------------------------------------------------------------------------
	output	 reg			Pulse;
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------
	//	State Encoding
	//--------------------------------------------------------------------------
	
	// place state encoding here
	
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Wire Declarations
	//--------------------------------------------------------------------------
	
	parameter INICIAL = 2'd00, INTERMEDIARIO = 2'd01, FINAL = 2'd11;

	// place wire declarations here	

	reg [1:0] state , proxState;
	
	always @(posedge Clock or negedge  Reset) begin

		if(!Reset) begin
			state <= INICIAL;
		end

		else state <= proxState;

	end

	always @(*) begin
		case(state)
		INICIAL:begin
			Pulse <= 0;
			if(Level == 0)begin
				proxState <= INTERMEDIARIO ;
			end
			else proxState <= INICIAL;
	
		end

		INTERMEDIARIO:begin
				Pulse <= 1;
				proxState <= FINAL;
		end

		FINAL:begin
			Pulse <= 1;
			if(Level == 1)begin
				proxState <= INICIAL ;
			end
			else proxState <= FINAL ;
		end

		endcase
	end


	//--------------------------------------------------------------------------
endmodule // LevelToPulse
module vga_controller(iRST_n,
                      iVGA_CLK,
							 codeColor,
                      oBLANK_n,
                      oHS,
                      oVS,
                      b_data,
                      g_data,
                      r_data);
input iRST_n;
input iVGA_CLK;
input [3:0] codeColor;
output reg oBLANK_n;
output reg oHS;
output reg oVS;
output [7:0] b_data;
output [7:0] g_data;  
output [7:0] r_data;                        
///////// ////                     
reg [18:0] ADDR;
reg [23:0] bgr_data;
wire VGA_CLK_n;
wire [7:0] index;
wire [23:0] bgr_data_raw;
wire cBLANK_n,cHS,cVS,rst;

reg [2:0]cor;
////
assign rst = ~iRST_n;
video_sync_generator LTM_ins (.vga_clk(iVGA_CLK),
                              .reset(rst),
                              .blank_n(cBLANK_n),
                              .HS(cHS),
                              .VS(cVS));
////
////Addresss generator
always@(posedge iVGA_CLK,negedge iRST_n)
begin
  if (!iRST_n)
     ADDR<=19'd0;
  else if (cHS==1'b0 && cVS==1'b0)
     ADDR<=19'd0;
  else if (cBLANK_n==1'b1)
     ADDR<=ADDR+1;
end
//////////////////////////
//////INDEX addr.
assign VGA_CLK_n = ~iVGA_CLK;
img_data	img_data_inst (
	.address ( ADDR ),
	.clock ( VGA_CLK_n ),
	.q ( index )
	);
//////Color table output
img_index	img_index_inst (
	.address ( index ),
	.clock ( iVGA_CLK ),
	.q ( bgr_data_raw)
	);	
//////
//////latch valid data at falling edge;
always@(posedge VGA_CLK_n) begin 

				bgr_data <= bgr_data_raw;
	
 			   if(bgr_data_raw == 24'he0) begin // Vermelho
					bgr_data <= 24'h0000AA;
				end 
				
				if(bgr_data_raw == 24'he0e0) begin  // Amarelog
					bgr_data <= 24'h00AAAA;
				end 
				
				if(bgr_data_raw == 24'hc04020) begin //Verde
					bgr_data <= 24'h007700;
				end
				
				if(bgr_data_raw == 24'h40a020) begin //Azul
					bgr_data <= 24'hAA0000;
				end 
				
				if(bgr_data_raw == 24'he0 && codeColor == 4'b0001 ) begin 
					bgr_data <= 24'h0000FF;
				end 
				
				if(bgr_data_raw == 24'he0e0 && codeColor == 4'b0011 ) begin 
					bgr_data <= 24'h00ffff;
				end
				
				if(bgr_data_raw == 24'hc04020 && codeColor == 4'b0010 ) begin 
					bgr_data <= 24'h00AA00;
				end
				
				if(bgr_data_raw == 24'h40a020 && codeColor == 4'b0100 ) begin 
					bgr_data <= 24'hff0000;
				end 
				
end 
assign b_data = bgr_data[23:16];
assign g_data = bgr_data[15:8];
assign r_data = bgr_data[7:0];
///////////////////
//////Delay the iHD, iVD,iDEN for one clock cycle;
always@(negedge iVGA_CLK)
begin
  oHS<=cHS;
  oVS<=cVS;
  oBLANK_n<=cBLANK_n;
end

endmodule
 	
















